//top_connection
//
//
//
//
//
`ifdef TX_CONNECT_RX

`endif

`ifdef PHY_BYPASS
`endif//`ifndef PHY_BYPASS

`ifdef MAC_BYPASS
`endif

`ifdef TX_SINGLE
`endif 

`ifdef RX_SINGLE
`endif

