//--------------------------------------------------------------------------
//interface
//--------------------------------------------------------------------------


`ifndef SUB_INTERFACE_SV
`define SUB_INTERFACE_SV

interface sub_interface #(parameter WIDTH = 8)(input bit = clk, input bit rst);
  logic pclk;
  assign pclk = clk;
  

endinterface

interface 
endinterface

interface    
endinterface


interface 
endinterface
  





`endif 
