`ifndef CONTROL_ENV
`define CONTROL_ENV



`endif 